module controller ();

endmodule
